// Defines the parameters for the system-level design

localparam PICASO_ID_WIDTH = 8;     // Row/Column ID width of PICASO blocks. 8bit: 256 x 256 x 16 PEs (2^20)
localparam NET_LEVEL_WIDTH = 3;     // width of net-level of PiCaSO's datanet-node
