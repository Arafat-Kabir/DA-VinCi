// defines the parameters of vvblock module
localparam VV_ACTCODE_WIDTH = 2;    // witdth of the activation table selection code
