// Defines the parameters for VV-Engine system-level design

localparam VVENG_RF_WIDTH = 16,
           VVENG_RF_DEPTH = 1024,
           VVENG_ID_WIDTH = 8;

